module webgpu

import webgpu.binding

pub struct Sampler {
	ptr binding.WGPUSampler
}