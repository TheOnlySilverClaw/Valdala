module binding

pub type WGPUQuerySet = voidptr

// TODO
