module binding

pub type WGPUComputePassEncoder = voidptr
pub type WGPUComputePipeline = voidptr

// TODO
