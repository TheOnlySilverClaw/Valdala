module binding