module binding

pub fn C.wgpuRenderPassEncoderEnd(encoder WGPURenderPassEncoder)

pub fn C.wgpuRenderPassEncoderRelease(encoder WGPURenderPassEncoder)
