module main

import log

import graphics


fn main() {

	graphics.create_renderer()!

	log.info("done")
}