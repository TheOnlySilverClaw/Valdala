module binding

#flag -I include

#include "wgpu.h"