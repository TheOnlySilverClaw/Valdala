module webgpu

#flag -L libraries

#flag -l c
#flag -l m
#flag -l wgpu_native
