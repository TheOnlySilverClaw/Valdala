module webgpu

// TODO