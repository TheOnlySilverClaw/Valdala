module webgpu

// TODO
