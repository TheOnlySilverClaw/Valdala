module binding

pub fn C.wgpuPipelineLayoutRelease(layout WGPUPipelineLayout)
