module webgpu

import webgpu.binding

pub struct Buffer {
	ptr binding.WGPUBuffer
}
