module binding

#flag -I include

#include "wgpu.h"

pub type WGPUBool = u32
