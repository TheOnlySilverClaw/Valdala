module webgpu

import webgpu.binding

pub struct PipelineLayout {
	ptr binding.WGPUPipelineLayout
}
