module binding
