module binding

// TODO
