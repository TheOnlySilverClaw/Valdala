module binding

pub fn C.wgpuCommandBufferRelease(buffer WGPUCommandBuffer)
