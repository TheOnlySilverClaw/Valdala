module binding

pub type WGPURenderBundle = voidptr
pub type WGPURenderBundleEncoder = voidptr

// TODO
