module binding

// TODO